
-- how colision works:
-- on vertical colision (colision with paddles) X velocity of the ball is inverted, Y velocity isnt changed
-- on horizontal colision (colision with top and botton of frame) X veloociity is constant, Y velocity is inverted

-- how are the clocks used:
-- pixel clock is used to output pixels of the ball
-- vsync is used to 

entity ball is  